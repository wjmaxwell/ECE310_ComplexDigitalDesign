// Test Bench for 3 Bit Full Adder

module fa3bit_tb;

  reg [2:0] A, B;
  wire [3:0] F;

  fa3bit DUT (
	A, B, F
  );

  initial begin
    $display( $time, ": A B | F" );
    $display( $time, ": ----+--" );
    $monitor( $time, ": %1d + %1d = %2d", A, B, F );
  end

  initial begin
        { A, B } = 6'b000_000;
    #10 { A, B } = 6'b000_001;
    #10 { A, B } = 6'b000_010;
    #10 { A, B } = 6'b000_011;
    #10 { A, B } = 6'b000_100;
    #10 { A, B } = 6'b000_101;
    #10 { A, B } = 6'b000_110;
    #10 { A, B } = 6'b000_111;

    #10 { A, B } = 6'b001_000;
    #10 { A, B } = 6'b001_001;
    #10 { A, B } = 6'b001_010;
    #10 { A, B } = 6'b001_011;
    #10 { A, B } = 6'b001_100;
    #10 { A, B } = 6'b001_101;
    #10 { A, B } = 6'b001_110;
    #10 { A, B } = 6'b001_111;

    #10 { A, B } = 6'b010_000;
    #10 { A, B } = 6'b010_001;
    #10 { A, B } = 6'b010_010;
    #10 { A, B } = 6'b010_011;
    #10 { A, B } = 6'b010_100;
    #10 { A, B } = 6'b010_101;
    #10 { A, B } = 6'b010_110;
    #10 { A, B } = 6'b010_111;

    #10 { A, B } = 6'b011_000;
    #10 { A, B } = 6'b011_001;
    #10 { A, B } = 6'b011_010;
    #10 { A, B } = 6'b011_011;
    #10 { A, B } = 6'b011_100;
    #10 { A, B } = 6'b011_101;
    #10 { A, B } = 6'b011_110;
    #10 { A, B } = 6'b011_111;

    #10 { A, B } = 6'b100_000;
    #10 { A, B } = 6'b100_001;
    #10 { A, B } = 6'b100_010;
    #10 { A, B } = 6'b100_011;
    #10 { A, B } = 6'b100_100;
    #10 { A, B } = 6'b100_101;
    #10 { A, B } = 6'b100_110;
    #10 { A, B } = 6'b100_111;

    #10 { A, B } = 6'b101_000;
    #10 { A, B } = 6'b101_001;
    #10 { A, B } = 6'b101_010;
    #10 { A, B } = 6'b101_011;
    #10 { A, B } = 6'b101_100;
    #10 { A, B } = 6'b101_101;
    #10 { A, B } = 6'b101_110;
    #10 { A, B } = 6'b101_111;

    #10 { A, B } = 6'b110_000;
    #10 { A, B } = 6'b110_001;
    #10 { A, B } = 6'b110_010;
    #10 { A, B } = 6'b110_011;
    #10 { A, B } = 6'b110_100;
    #10 { A, B } = 6'b110_101;
    #10 { A, B } = 6'b110_110;
    #10 { A, B } = 6'b110_111;

    #10 { A, B } = 6'b111_000;
    #10 { A, B } = 6'b111_001;
    #10 { A, B } = 6'b111_010;
    #10 { A, B } = 6'b111_011;
    #10 { A, B } = 6'b111_100;
    #10 { A, B } = 6'b111_101;
    #10 { A, B } = 6'b111_110;
    #10 { A, B } = 6'b111_111;

    #10 $stop();
  end

endmodule
